module and_gate(A,B,Y);
input A,B;
output Y;
    and(Y, A, B);
endmodule
